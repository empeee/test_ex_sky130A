magic
tech sky130A
timestamp 1747405320
<< locali >>
rect 112 1084 384 1116
rect -48 -50 48 98
rect 528 -50 624 98
rect -100 -55 650 -50
rect -100 -145 147 -55
rect 237 -145 650 -55
rect -100 -150 650 -145
<< viali >>
rect 147 -145 237 -55
<< metal1 >>
rect 500 1912 600 2000
rect 336 1816 600 1912
rect 80 1116 112 1716
rect 77 1084 80 1116
rect 112 1084 115 1116
rect 80 284 112 1084
rect 144 -55 240 1798
rect 500 1512 600 1816
rect 336 1416 600 1512
rect 384 1116 416 1119
rect 384 1081 416 1084
rect 500 748 600 1416
rect 336 652 600 748
rect 500 348 600 652
rect 336 252 600 348
rect 500 0 600 252
rect 144 -145 147 -55
rect 237 -145 240 -55
rect 144 -151 240 -145
<< via1 >>
rect 80 1084 112 1116
rect 384 1084 416 1116
<< metal2 >>
rect 80 1116 112 1119
rect 112 1084 384 1116
rect 416 1084 419 1116
rect 80 1081 112 1084
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1740610800
transform 1 0 0 0 1 400
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1740610800
transform 1 0 0 0 1 1200
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1740610800
transform 1 0 0 0 1 800
box -92 -64 668 464
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1740610800
transform 1 0 0 0 1 1600
box -92 -64 668 464
<< labels >>
flabel locali -100 -150 650 -50 0 FreeSans 800 0 0 0 VSS
flabel metal1 336 1816 600 1912 0 FreeSans 800 0 0 0 IBNS_20U
port 2 nsew
flabel metal2 112 1084 384 1116 0 FreeSans 800 0 0 0 IBPS_5U
port 4 nsew
flabel locali 237 -150 650 -50 0 FreeSans 800 0 0 0 VSS
port 6 nsew
<< end >>
